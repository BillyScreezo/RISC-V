/***********************************************************************************
 * Copyright (C) 2024 Kirill Turintsev <billiscreezo228@gmail.com>
 * See LICENSE file for licensing details.
 *
 * This file contains declarations for the INTCTRL module
 *
 ***********************************************************************************/
 
 package riscv_intc_pkg;
	
	parameter int NUMINT = 4;

endpackage : riscv_intc_pkg